`timescale 1ns / 1ps

module mem_reader_tb;

    axi_reader_v1_0 uut (
        
    );

endmodule
